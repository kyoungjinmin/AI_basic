library verilog;
use verilog.vl_types.all;
entity tb_hw_assign is
end tb_hw_assign;
