library verilog;
use verilog.vl_types.all;
entity pencase_seq_tb is
end pencase_seq_tb;
