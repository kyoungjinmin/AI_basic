library verilog;
use verilog.vl_types.all;
entity doorlock_2_tb is
end doorlock_2_tb;
