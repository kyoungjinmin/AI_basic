library verilog;
use verilog.vl_types.all;
entity practice_tb is
end practice_tb;
