library verilog;
use verilog.vl_types.all;
entity doorlock_tb is
end doorlock_tb;
