library verilog;
use verilog.vl_types.all;
entity always_tb is
end always_tb;
