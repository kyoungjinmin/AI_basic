library verilog;
use verilog.vl_types.all;
entity tb_final_123 is
end tb_final_123;
