library verilog;
use verilog.vl_types.all;
entity tb_hw is
end tb_hw;
