library verilog;
use verilog.vl_types.all;
entity tb_final_359 is
end tb_final_359;
